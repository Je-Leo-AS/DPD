--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_textio.ALL;
USE std.textio.ALL;

ENTITY tb IS
END tb;
 
ARCHITECTURE behavior OF tb IS 
    CONSTANT n_bits_resolution : INTEGER := 9;
    CONSTANT n_bits_overflow : INTEGER := 8;
    CONSTANT n_signals_used : INTEGER := 2;
    CONSTANT n_polygnos_degree : INTEGER := 2;
    -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT dpd
        PORT (
            reset : IN STD_LOGIC;
            clk : IN STD_LOGIC;
            UR : IN STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);
            UI : IN STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);
            UR_out : OUT STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);
            UI_out : OUT STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0)
        );
    END COMPONENT;

    -- Signals for connecting to UUT
    SIGNAL reset : STD_LOGIC := '0';
    SIGNAL clk : STD_LOGIC := '0';
    SIGNAL UR : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL UI : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL UR_out : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL UI_out : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);

    -- Clock period definition
    CONSTANT clk_period : TIME := 16 ns;
    FILE output_file : TEXT OPEN WRITE_MODE IS "simulation_output.txt";
    SHARED VARIABLE line_buffer : LINE;
    SHARED VARIABLE data : INTEGER;

 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: DPD PORT MAP (
          reset => reset,
          clk => clk,
          UR => UR,
          UI => UI,
          UR_out => UR_out,
          UI_out => UI_out
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   write_output : PROCESS
   BEGIN
      IF reset = '1' THEN
		
    ELSIF rising_edge(clk) THEN
        WRITE(line_buffer, to_integer(UR_out));
        WRITE(line_buffer, STRING'(" + "));
        WRITE(line_buffer, to_integer(UI_out));
        WRITE(line_buffer, STRING'("j"));
        WRITELINE(output_file, line_buffer);
    END IF;
   END PROCESS;

      -- in process
   calc_proc: process
   begin		
      reset <= '1';
      wait for 2 * clk_period;	
      reset <= '0';
      WAIT FOR clk_period;
      
UR <= "000111101";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "010100001";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "010001000";
WAIT FOR clk_period;
UR <= "110100101";
UI <= "001110100";
WAIT FOR clk_period;
UR <= "110001111";
UI <= "001011110";
WAIT FOR clk_period;
UR <= "101111110";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000011100";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000101111";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "101100010";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000111111";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "101010000";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "101001011";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "101000111";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "101001001";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000011000";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "110000011";
UI <= "001010000";
WAIT FOR clk_period;
UR <= "110011110";
UI <= "001110010";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "010010011";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "111111000";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "011001011";
WAIT FOR clk_period;
UR <= "000101000";
UI <= "011000011";
WAIT FOR clk_period;
UR <= "000111000";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "010000111";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "001010101";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "110101101";
WAIT FOR clk_period;
UR <= "000000110";
UI <= "110000000";
WAIT FOR clk_period;
UR <= "111101111";
UI <= "101011100";
WAIT FOR clk_period;
UR <= "111010110";
UI <= "101001010";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "110001111";
UI <= "101110001";
WAIT FOR clk_period;
UR <= "101111101";
UI <= "110010110";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "111000001";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "000010000";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "000101111";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "001000101";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "110000011";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "110010100";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "111100011";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "111001010";
UI <= "110001101";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "101100110";
WAIT FOR clk_period;
UR <= "111011110";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "111100100";
UI <= "100101001";
WAIT FOR clk_period;
UR <= "111100011";
UI <= "100011000";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "100010000";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "100001111";
WAIT FOR clk_period;
UR <= "111010011";
UI <= "100011010";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "100101011";
WAIT FOR clk_period;
UR <= "111000110";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "111000111";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "110000001";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "111100101";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "111110110";
UI <= "111110100";
WAIT FOR clk_period;
UR <= "000001010";
UI <= "000011011";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "001100101";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "000111001";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "011010001";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "011010100";
WAIT FOR clk_period;
UR <= "000010001";
UI <= "011010001";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "011001001";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "010111100";
WAIT FOR clk_period;
UR <= "000001001";
UI <= "010101011";
WAIT FOR clk_period;
UR <= "000010111";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "000101110";
UI <= "010000001";
WAIT FOR clk_period;
UR <= "001001110";
UI <= "001101010";
WAIT FOR clk_period;
UR <= "001101111";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "010010010";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "010110000";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "011000011";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "011001011";
UI <= "111110100";
WAIT FOR clk_period;
UR <= "011000101";
UI <= "111011111";
WAIT FOR clk_period;
UR <= "010110000";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "110110010";
WAIT FOR clk_period;
UR <= "001100100";
UI <= "110011100";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "110001010";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "101111011";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "101100100";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "101011100";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "101011100";
WAIT FOR clk_period;
UR <= "111000111";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "111101001";
UI <= "101101000";
WAIT FOR clk_period;
UR <= "000010111";
UI <= "101110011";
WAIT FOR clk_period;
UR <= "001001001";
UI <= "110000011";
WAIT FOR clk_period;
UR <= "001111001";
UI <= "110010100";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "110100110";
WAIT FOR clk_period;
UR <= "010111110";
UI <= "110111100";
WAIT FOR clk_period;
UR <= "011001000";
UI <= "111001110";
WAIT FOR clk_period;
UR <= "010111100";
UI <= "111011110";
WAIT FOR clk_period;
UR <= "010011111";
UI <= "111101111";
WAIT FOR clk_period;
UR <= "001110000";
UI <= "111111110";
WAIT FOR clk_period;
UR <= "000110111";
UI <= "000001001";
WAIT FOR clk_period;
UR <= "111110110";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101011000";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101000000";
UI <= "000101000";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "000101000";
WAIT FOR clk_period;
UR <= "101111011";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "000011101";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "000101100";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "001101001";
UI <= "111111110";
WAIT FOR clk_period;
UR <= "010011010";
UI <= "111101101";
WAIT FOR clk_period;
UR <= "010111111";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "011010000";
UI <= "111000010";
WAIT FOR clk_period;
UR <= "011010000";
UI <= "110101100";
WAIT FOR clk_period;
UR <= "010111111";
UI <= "110010110";
WAIT FOR clk_period;
UR <= "010011101";
UI <= "110000000";
WAIT FOR clk_period;
UR <= "001110010";
UI <= "101101110";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "000001101";
UI <= "101010110";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "110101110";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "110001011";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "101111010";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "110010011";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "110110010";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "111010010";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "111110010";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000010001";
WAIT FOR clk_period;
UR <= "101101100";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101111100";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "110001010";
UI <= "001011011";
WAIT FOR clk_period;
UR <= "110011010";
UI <= "001101001";
WAIT FOR clk_period;
UR <= "110101100";
UI <= "001110100";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "111010100";
UI <= "010000001";
WAIT FOR clk_period;
UR <= "111101010";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "010001010";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010010000";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "001001101";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "001011111";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "001101010";
UI <= "010111011";
WAIT FOR clk_period;
UR <= "001101110";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "011001001";
WAIT FOR clk_period;
UR <= "001011110";
UI <= "011001000";
WAIT FOR clk_period;
UR <= "001000111";
UI <= "010111111";
WAIT FOR clk_period;
UR <= "000101011";
UI <= "010110000";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "010011001";
WAIT FOR clk_period;
UR <= "111100100";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "110111110";
UI <= "001011110";
WAIT FOR clk_period;
UR <= "110011101";
UI <= "001000010";
WAIT FOR clk_period;
UR <= "110000000";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "101101001";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000001111";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "101101110";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "110000100";
UI <= "001010101";
WAIT FOR clk_period;
UR <= "110011111";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "110111110";
UI <= "010011011";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "111111011";
UI <= "011001000";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "011001100";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "010111110";
WAIT FOR clk_period;
UR <= "000111010";
UI <= "010100010";
WAIT FOR clk_period;
UR <= "001000010";
UI <= "001110110";
WAIT FOR clk_period;
UR <= "001000101";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "000111111";
UI <= "000000110";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "000100001";
UI <= "110010010";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "101001011";
WAIT FOR clk_period;
UR <= "111010000";
UI <= "101000001";
WAIT FOR clk_period;
UR <= "110110010";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "110010101";
UI <= "101100001";
WAIT FOR clk_period;
UR <= "101111011";
UI <= "110000110";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "110110011";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "111100010";
WAIT FOR clk_period;
UR <= "101001110";
UI <= "000001110";
WAIT FOR clk_period;
UR <= "101001101";
UI <= "000110000";
WAIT FOR clk_period;

      -- insert stimulus here 
      wait;
   end process;
    
END;
