--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE ieee.std_logic_textio.ALL;
USE std.textio.ALL;
LIBRARY work;
USE work.functions_Package.ALL;

ENTITY tb IS
END tb;
 
ARCHITECTURE behavior OF tb IS 
    -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT dpd
        PORT (
            reset : IN STD_LOGIC;
            clk : IN STD_LOGIC;
            UR : IN STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);
            UI : IN STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);
            UR_out : OUT STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);
            UI_out : OUT STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0)
        );
    END COMPONENT;

    -- Signals for connecting to UUT
    SIGNAL reset : STD_LOGIC := '0';
    SIGNAL clk : STD_LOGIC := '0';
    SIGNAL UR : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL UI : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL UR_out : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL UI_out : STD_LOGIC_VECTOR(n_bits_resolution - 1 DOWNTO 0);

    -- Clock period definition
    CONSTANT clk_period : TIME := 16 ns;
    FILE output_file : TEXT OPEN WRITE_MODE IS "simulation_output.txt";
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: DPD PORT MAP (
          reset => reset,
          clk => clk,
          UR => UR,
          UI => UI,
          UR_out => UR_out,
          UI_out => UI_out
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
    write_output : PROCESS(clk)
        VARIABLE line_buffer : LINE;
        VARIABLE data : INTEGER;
    BEGIN
        IF reset = '0' and rising_edge(clk) THEN
            WRITE(line_buffer, to_integer(signed(UR_out)));
            WRITE(line_buffer, STRING'(","));
            WRITE(line_buffer, to_integer(signed(UI_out)));
            WRITE(line_buffer, STRING'("j"));
            WRITELINE(output_file, line_buffer);
        END IF;
    END PROCESS;

      -- in process
   calc_proc: process
   begin		
      reset <= '1';
      wait for 2 * clk_period;	
      reset <= '0';
      WAIT FOR clk_period;
      
UR <= "000111101";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "010100001";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "010001000";
WAIT FOR clk_period;
UR <= "110100101";
UI <= "001110100";
WAIT FOR clk_period;
UR <= "110001111";
UI <= "001011110";
WAIT FOR clk_period;
UR <= "101111110";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000011100";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000101111";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "101100010";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000111111";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "101010000";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "101001011";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "101000111";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "101001001";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000011000";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "110000011";
UI <= "001010000";
WAIT FOR clk_period;
UR <= "110011110";
UI <= "001110010";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "010010011";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "111111000";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "011001011";
WAIT FOR clk_period;
UR <= "000101000";
UI <= "011000011";
WAIT FOR clk_period;
UR <= "000111000";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "010000111";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "001010101";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "110101101";
WAIT FOR clk_period;
UR <= "000000110";
UI <= "110000000";
WAIT FOR clk_period;
UR <= "111101111";
UI <= "101011100";
WAIT FOR clk_period;
UR <= "111010110";
UI <= "101001010";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "110001111";
UI <= "101110001";
WAIT FOR clk_period;
UR <= "101111101";
UI <= "110010110";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "111000001";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "000010000";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "000101111";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "001000101";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "110000011";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "110010100";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "111100011";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "111001010";
UI <= "110001101";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "101100110";
WAIT FOR clk_period;
UR <= "111011110";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "111100100";
UI <= "100101001";
WAIT FOR clk_period;
UR <= "111100011";
UI <= "100011000";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "100010000";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "100001111";
WAIT FOR clk_period;
UR <= "111010011";
UI <= "100011010";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "100101011";
WAIT FOR clk_period;
UR <= "111000110";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "111000111";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "110000001";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "111100101";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "111110110";
UI <= "111110100";
WAIT FOR clk_period;
UR <= "000001010";
UI <= "000011011";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "001100101";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "000111001";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "011010001";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "011010100";
WAIT FOR clk_period;
UR <= "000010001";
UI <= "011010001";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "011001001";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "010111100";
WAIT FOR clk_period;
UR <= "000001001";
UI <= "010101011";
WAIT FOR clk_period;
UR <= "000010111";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "000101110";
UI <= "010000001";
WAIT FOR clk_period;
UR <= "001001110";
UI <= "001101010";
WAIT FOR clk_period;
UR <= "001101111";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "010010010";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "010110000";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "011000011";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "011001011";
UI <= "111110100";
WAIT FOR clk_period;
UR <= "011000101";
UI <= "111011111";
WAIT FOR clk_period;
UR <= "010110000";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "110110010";
WAIT FOR clk_period;
UR <= "001100100";
UI <= "110011100";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "110001010";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "101111011";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "101100100";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "101011100";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "101011100";
WAIT FOR clk_period;
UR <= "111000111";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "111101001";
UI <= "101101000";
WAIT FOR clk_period;
UR <= "000010111";
UI <= "101110011";
WAIT FOR clk_period;
UR <= "001001001";
UI <= "110000011";
WAIT FOR clk_period;
UR <= "001111001";
UI <= "110010100";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "110100110";
WAIT FOR clk_period;
UR <= "010111110";
UI <= "110111100";
WAIT FOR clk_period;
UR <= "011001000";
UI <= "111001110";
WAIT FOR clk_period;
UR <= "010111100";
UI <= "111011110";
WAIT FOR clk_period;
UR <= "010011111";
UI <= "111101111";
WAIT FOR clk_period;
UR <= "001110000";
UI <= "111111110";
WAIT FOR clk_period;
UR <= "000110111";
UI <= "000001001";
WAIT FOR clk_period;
UR <= "111110110";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101011000";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101000000";
UI <= "000101000";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "000101000";
WAIT FOR clk_period;
UR <= "101111011";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "000011101";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "000101100";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "001101001";
UI <= "111111110";
WAIT FOR clk_period;
UR <= "010011010";
UI <= "111101101";
WAIT FOR clk_period;
UR <= "010111111";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "011010000";
UI <= "111000010";
WAIT FOR clk_period;
UR <= "011010000";
UI <= "110101100";
WAIT FOR clk_period;
UR <= "010111111";
UI <= "110010110";
WAIT FOR clk_period;
UR <= "010011101";
UI <= "110000000";
WAIT FOR clk_period;
UR <= "001110010";
UI <= "101101110";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "000001101";
UI <= "101010110";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "110101110";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "110001011";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "101111010";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "110010011";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "110110010";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "111010010";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "111110010";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000010001";
WAIT FOR clk_period;
UR <= "101101100";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101111100";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "110001010";
UI <= "001011011";
WAIT FOR clk_period;
UR <= "110011010";
UI <= "001101001";
WAIT FOR clk_period;
UR <= "110101100";
UI <= "001110100";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "111010100";
UI <= "010000001";
WAIT FOR clk_period;
UR <= "111101010";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "010001010";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010010000";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "001001101";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "001011111";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "001101010";
UI <= "010111011";
WAIT FOR clk_period;
UR <= "001101110";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "011001001";
WAIT FOR clk_period;
UR <= "001011110";
UI <= "011001000";
WAIT FOR clk_period;
UR <= "001000111";
UI <= "010111111";
WAIT FOR clk_period;
UR <= "000101011";
UI <= "010110000";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "010011001";
WAIT FOR clk_period;
UR <= "111100100";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "110111110";
UI <= "001011110";
WAIT FOR clk_period;
UR <= "110011101";
UI <= "001000010";
WAIT FOR clk_period;
UR <= "110000000";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "101101001";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000001111";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "101101110";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "110000100";
UI <= "001010101";
WAIT FOR clk_period;
UR <= "110011111";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "110111110";
UI <= "010011011";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "111111011";
UI <= "011001000";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "011001100";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "010111110";
WAIT FOR clk_period;
UR <= "000111010";
UI <= "010100010";
WAIT FOR clk_period;
UR <= "001000010";
UI <= "001110110";
WAIT FOR clk_period;
UR <= "001000101";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "000111111";
UI <= "000000110";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "000100001";
UI <= "110010010";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "101001011";
WAIT FOR clk_period;
UR <= "111010000";
UI <= "101000001";
WAIT FOR clk_period;
UR <= "110110010";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "110010101";
UI <= "101100001";
WAIT FOR clk_period;
UR <= "101111011";
UI <= "110000110";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "110110011";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "111100010";
WAIT FOR clk_period;
UR <= "101001110";
UI <= "000001110";
WAIT FOR clk_period;
UR <= "101001101";
UI <= "000110000";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "001000101";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "001001011";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "110001010";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "110100001";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "110111001";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "111001010";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "101111100";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "111011111";
UI <= "101000101";
WAIT FOR clk_period;
UR <= "111010111";
UI <= "100111110";
WAIT FOR clk_period;
UR <= "111000101";
UI <= "101000110";
WAIT FOR clk_period;
UR <= "110110000";
UI <= "101011011";
WAIT FOR clk_period;
UR <= "110011010";
UI <= "101111101";
WAIT FOR clk_period;
UR <= "110000010";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "101101011";
UI <= "111010011";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "001001011";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "001100101";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "001110110";
WAIT FOR clk_period;
UR <= "110001110";
UI <= "010000001";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "111110011";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "010000110";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "010001001";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "010001110";
WAIT FOR clk_period;
UR <= "001001100";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "001001111";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "001001100";
UI <= "010110010";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "010111110";
WAIT FOR clk_period;
UR <= "000111000";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "011001001";
WAIT FOR clk_period;
UR <= "000100100";
UI <= "011000010";
WAIT FOR clk_period;
UR <= "000011111";
UI <= "010110101";
WAIT FOR clk_period;
UR <= "000011111";
UI <= "010100001";
WAIT FOR clk_period;
UR <= "000100110";
UI <= "010000100";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "001100011";
WAIT FOR clk_period;
UR <= "001000101";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "001011011";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "001110011";
UI <= "111111111";
WAIT FOR clk_period;
UR <= "010001010";
UI <= "111100011";
WAIT FOR clk_period;
UR <= "010100000";
UI <= "111001111";
WAIT FOR clk_period;
UR <= "010110010";
UI <= "111000100";
WAIT FOR clk_period;
UR <= "010111110";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "011000101";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "011000101";
UI <= "111001010";
WAIT FOR clk_period;
UR <= "011000010";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "010111011";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "010110010";
UI <= "111101001";
WAIT FOR clk_period;
UR <= "010100101";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "010011001";
UI <= "111101000";
WAIT FOR clk_period;
UR <= "010001101";
UI <= "111011111";
WAIT FOR clk_period;
UR <= "001111111";
UI <= "111001101";
WAIT FOR clk_period;
UR <= "001110010";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "001100101";
UI <= "110011110";
WAIT FOR clk_period;
UR <= "001010100";
UI <= "110000101";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "000101000";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "000001100";
UI <= "101010000";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "101001110";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "101011000";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "101101011";
WAIT FOR clk_period;
UR <= "101111110";
UI <= "110000101";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "101000110";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "100110101";
UI <= "111110001";
WAIT FOR clk_period;
UR <= "100110001";
UI <= "000010010";
WAIT FOR clk_period;
UR <= "100111011";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000111111";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "001001001";
WAIT FOR clk_period;
UR <= "110100001";
UI <= "001000111";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "000001011";
UI <= "000101100";
WAIT FOR clk_period;
UR <= "000111111";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "001110000";
UI <= "111111010";
WAIT FOR clk_period;
UR <= "010010100";
UI <= "111100010";
WAIT FOR clk_period;
UR <= "010101100";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "010110111";
UI <= "110111001";
WAIT FOR clk_period;
UR <= "010110011";
UI <= "110101010";
WAIT FOR clk_period;
UR <= "010011111";
UI <= "110100001";
WAIT FOR clk_period;
UR <= "010000001";
UI <= "110011101";
WAIT FOR clk_period;
UR <= "001011011";
UI <= "110011000";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "110010101";
WAIT FOR clk_period;
UR <= "000001011";
UI <= "110001111";
WAIT FOR clk_period;
UR <= "111100111";
UI <= "110000101";
WAIT FOR clk_period;
UR <= "111001000";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "101010010";
WAIT FOR clk_period;
UR <= "110100101";
UI <= "101000000";
WAIT FOR clk_period;
UR <= "110101010";
UI <= "100101101";
WAIT FOR clk_period;
UR <= "110110101";
UI <= "100100000";
WAIT FOR clk_period;
UR <= "111000010";
UI <= "100011100";
WAIT FOR clk_period;
UR <= "111010001";
UI <= "100100001";
WAIT FOR clk_period;
UR <= "111011110";
UI <= "100110001";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "101001111";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "101110111";
WAIT FOR clk_period;
UR <= "111110000";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "111110000";
UI <= "111011101";
WAIT FOR clk_period;
UR <= "111110001";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "111110100";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "111111000";
UI <= "001110101";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "000010010";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "000101001";
UI <= "010110010";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "010101010";
WAIT FOR clk_period;
UR <= "001011100";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "001110101";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "001010100";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "010101110";
UI <= "000001010";
WAIT FOR clk_period;
UR <= "010110001";
UI <= "111101001";
WAIT FOR clk_period;
UR <= "010101010";
UI <= "111010000";
WAIT FOR clk_period;
UR <= "010011010";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "010000000";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "001011111";
UI <= "110111010";
WAIT FOR clk_period;
UR <= "000111000";
UI <= "111000101";
WAIT FOR clk_period;
UR <= "000001100";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "111101011";
WAIT FOR clk_period;
UR <= "110110100";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "110001001";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000110000";
WAIT FOR clk_period;
UR <= "101000000";
UI <= "001000011";
WAIT FOR clk_period;
UR <= "100100011";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "100001111";
UI <= "001011100";
WAIT FOR clk_period;
UR <= "100000011";
UI <= "001100001";
WAIT FOR clk_period;
UR <= "100000000";
UI <= "001100001";
WAIT FOR clk_period;
UR <= "100001010";
UI <= "001011010";
WAIT FOR clk_period;
UR <= "100011100";
UI <= "001001101";
WAIT FOR clk_period;
UR <= "100111010";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "110010000";
UI <= "000010010";
WAIT FOR clk_period;
UR <= "111000101";
UI <= "111111010";
WAIT FOR clk_period;
UR <= "111111100";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "111001110";
WAIT FOR clk_period;
UR <= "001100010";
UI <= "111000001";
WAIT FOR clk_period;
UR <= "010001010";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "010100111";
UI <= "110111001";
WAIT FOR clk_period;
UR <= "010110101";
UI <= "111000010";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "010101001";
UI <= "111110010";
WAIT FOR clk_period;
UR <= "010010010";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "001110011";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "001010100";
UI <= "001100001";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "010000100";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "000001111";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "000001110";
UI <= "010110101";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "001010011";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "001111010";
UI <= "001010001";
WAIT FOR clk_period;
UR <= "010011110";
UI <= "000101010";
WAIT FOR clk_period;
UR <= "010111010";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "011001010";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "011001010";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "010111010";
UI <= "110111010";
WAIT FOR clk_period;
UR <= "010011000";
UI <= "110111001";
WAIT FOR clk_period;
UR <= "001101000";
UI <= "111000100";
WAIT FOR clk_period;
UR <= "000101011";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "111110001";
WAIT FOR clk_period;
UR <= "110110000";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "101111011";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "101000001";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "101010111";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "101111111";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "110110100";
UI <= "000001110";
WAIT FOR clk_period;
UR <= "111110011";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "000110000";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "001101010";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "010011011";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "010111110";
UI <= "110111100";
WAIT FOR clk_period;
UR <= "011001110";
UI <= "111001010";
WAIT FOR clk_period;
UR <= "011001111";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "011000000";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "010000100";
UI <= "001010011";
WAIT FOR clk_period;
UR <= "001011111";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "000111101";
UI <= "010011000";
WAIT FOR clk_period;
UR <= "000100000";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "000001110";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "010110100";
WAIT FOR clk_period;
UR <= "000001101";
UI <= "010100011";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "010001001";
WAIT FOR clk_period;
UR <= "000110110";
UI <= "001100111";
WAIT FOR clk_period;
UR <= "001010100";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "001110100";
UI <= "000011001";
WAIT FOR clk_period;
UR <= "010010100";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "010101111";
UI <= "111010010";
WAIT FOR clk_period;
UR <= "011000011";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "011001111";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "011010011";
UI <= "110011010";
WAIT FOR clk_period;
UR <= "011010000";
UI <= "110011000";
WAIT FOR clk_period;
UR <= "011001000";
UI <= "110011101";
WAIT FOR clk_period;
UR <= "010111011";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "010101011";
UI <= "110110110";
WAIT FOR clk_period;
UR <= "010011101";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "010010000";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "010000010";
UI <= "111110001";
WAIT FOR clk_period;
UR <= "001111010";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "001110001";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "000110111";
WAIT FOR clk_period;
UR <= "001100101";
UI <= "001001101";
WAIT FOR clk_period;
UR <= "001011100";
UI <= "001100101";
WAIT FOR clk_period;
UR <= "001010100";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "001001000";
UI <= "010010000";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "010100100";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "010110011";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "010111101";
WAIT FOR clk_period;
UR <= "000001010";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "111111110";
UI <= "011000111";
WAIT FOR clk_period;
UR <= "111111000";
UI <= "011000100";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "010111110";
WAIT FOR clk_period;
UR <= "000000000";
UI <= "010110010";
WAIT FOR clk_period;
UR <= "000010000";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "000100110";
UI <= "010010100";
WAIT FOR clk_period;
UR <= "001000010";
UI <= "010000000";
WAIT FOR clk_period;
UR <= "001100100";
UI <= "001101101";
WAIT FOR clk_period;
UR <= "010000100";
UI <= "001011000";
WAIT FOR clk_period;
UR <= "010100001";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "011000100";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "011000100";
UI <= "111111100";
WAIT FOR clk_period;
UR <= "010111001";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "010100001";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "001111111";
UI <= "110101010";
WAIT FOR clk_period;
UR <= "001011000";
UI <= "110010000";
WAIT FOR clk_period;
UR <= "000101100";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "000000011";
UI <= "101100100";
WAIT FOR clk_period;
UR <= "111100010";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "101001100";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "101001110";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "111001111";
UI <= "101100100";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "000010010";
UI <= "110010001";
WAIT FOR clk_period;
UR <= "000111110";
UI <= "110101001";
WAIT FOR clk_period;
UR <= "001101001";
UI <= "111000000";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "010101011";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "010111000";
UI <= "111100101";
WAIT FOR clk_period;
UR <= "010111000";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "010101000";
UI <= "111010011";
WAIT FOR clk_period;
UR <= "010001100";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "001100100";
UI <= "110101000";
WAIT FOR clk_period;
UR <= "000111001";
UI <= "110001101";
WAIT FOR clk_period;
UR <= "000010000";
UI <= "101110100";
WAIT FOR clk_period;
UR <= "111101000";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "111001100";
UI <= "101010010";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "101001101";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "101010010";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "111100111";
UI <= "101110101";
WAIT FOR clk_period;
UR <= "000001100";
UI <= "110010001";
WAIT FOR clk_period;
UR <= "000110110";
UI <= "110101100";
WAIT FOR clk_period;
UR <= "001100001";
UI <= "111000101";
WAIT FOR clk_period;
UR <= "010001001";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "010101001";
UI <= "111100101";
WAIT FOR clk_period;
UR <= "010111010";
UI <= "111101000";
WAIT FOR clk_period;
UR <= "011000000";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "010110101";
UI <= "111010001";
WAIT FOR clk_period;
UR <= "010011111";
UI <= "110111001";
WAIT FOR clk_period;
UR <= "001111110";
UI <= "110011101";
WAIT FOR clk_period;
UR <= "001010101";
UI <= "110000010";
WAIT FOR clk_period;
UR <= "000100111";
UI <= "101101000";
WAIT FOR clk_period;
UR <= "111111101";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "111010011";
UI <= "101001100";
WAIT FOR clk_period;
UR <= "110110000";
UI <= "101001100";
WAIT FOR clk_period;
UR <= "110010100";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "101110001";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "110010000";
WAIT FOR clk_period;
UR <= "101101110";
UI <= "110110101";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "101110001";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101110001";
UI <= "000111100";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "001001110";
WAIT FOR clk_period;
UR <= "101101110";
UI <= "001010110";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "001010110";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "001001111";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "001000010";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "101010000";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000011111";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000011000";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101110010";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "000111100";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "000111111";
WAIT FOR clk_period;
UR <= "101100101";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101000100";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "100111100";
UI <= "000001111";
WAIT FOR clk_period;
UR <= "100110111";
UI <= "000000111";
WAIT FOR clk_period;
UR <= "100111010";
UI <= "000000110";
WAIT FOR clk_period;
UR <= "101000001";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000011000";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "110100000";
UI <= "001100010";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "001111110";
WAIT FOR clk_period;
UR <= "111100001";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "111111110";
UI <= "010101010";
WAIT FOR clk_period;
UR <= "000010110";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "000101000";
UI <= "010111000";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "010101011";
WAIT FOR clk_period;
UR <= "000110110";
UI <= "010010101";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "001110100";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "000011011";
WAIT FOR clk_period;
UR <= "000001100";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "110111110";
WAIT FOR clk_period;
UR <= "111100111";
UI <= "110010000";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "101101011";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "101001110";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "100111000";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "100101100";
WAIT FOR clk_period;
UR <= "110111011";
UI <= "100101000";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "100101101";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "100110100";
WAIT FOR clk_period;
UR <= "111001000";
UI <= "101000000";
WAIT FOR clk_period;
UR <= "111001110";
UI <= "101010001";
WAIT FOR clk_period;
UR <= "111010100";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "111011111";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "111100010";
UI <= "110000000";
WAIT FOR clk_period;
UR <= "111100101";
UI <= "110000100";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "110000100";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "101111110";
WAIT FOR clk_period;
UR <= "111100010";
UI <= "101110110";
WAIT FOR clk_period;
UR <= "111011110";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "111010001";
UI <= "101010000";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "111000011";
UI <= "100111000";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "100101111";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "100101101";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "100110000";
WAIT FOR clk_period;
UR <= "110111010";
UI <= "100111010";
WAIT FOR clk_period;
UR <= "111000010";
UI <= "101001100";
WAIT FOR clk_period;
UR <= "111001111";
UI <= "101100110";
WAIT FOR clk_period;
UR <= "111100001";
UI <= "110000111";
WAIT FOR clk_period;
UR <= "111110101";
UI <= "110101101";
WAIT FOR clk_period;
UR <= "000001011";
UI <= "111011000";
WAIT FOR clk_period;
UR <= "000100000";
UI <= "000000110";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "000111110";
UI <= "001011101";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "010000001";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "010011111";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "010110100";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "010111101";
WAIT FOR clk_period;
UR <= "111111100";
UI <= "010111101";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "010110010";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "110001100";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "101101010";
UI <= "001100110";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "101001000";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "101001000";
UI <= "000000100";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "111100101";
WAIT FOR clk_period;
UR <= "101100111";
UI <= "111001010";
WAIT FOR clk_period;
UR <= "110000100";
UI <= "110110011";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "110011111";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "110001110";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "101111111";
WAIT FOR clk_period;
UR <= "111101010";
UI <= "101110011";
WAIT FOR clk_period;
UR <= "111110010";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "111110000";
UI <= "101011011";
WAIT FOR clk_period;
UR <= "111100101";
UI <= "101010010";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "110110000";
UI <= "101000000";
WAIT FOR clk_period;
UR <= "110100100";
UI <= "101000010";
WAIT FOR clk_period;
UR <= "110100010";
UI <= "101000111";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "101010001";
WAIT FOR clk_period;
UR <= "111000110";
UI <= "101011110";
WAIT FOR clk_period;
UR <= "111101001";
UI <= "101101111";
WAIT FOR clk_period;
UR <= "000010010";
UI <= "110000011";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "110010101";
WAIT FOR clk_period;
UR <= "001110011";
UI <= "110101001";
WAIT FOR clk_period;
UR <= "010011011";
UI <= "110111011";
WAIT FOR clk_period;
UR <= "010111000";
UI <= "111001001";
WAIT FOR clk_period;
UR <= "011000101";
UI <= "111010100";
WAIT FOR clk_period;
UR <= "011000010";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "010101010";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "010000011";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "001010000";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "000010101";
UI <= "111101001";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "111110000";
WAIT FOR clk_period;
UR <= "110100010";
UI <= "111111001";
WAIT FOR clk_period;
UR <= "101110010";
UI <= "000000110";
WAIT FOR clk_period;
UR <= "101010010";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101000011";
UI <= "000101100";
WAIT FOR clk_period;
UR <= "101000011";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "001011110";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "001110110";
WAIT FOR clk_period;
UR <= "110011010";
UI <= "010001101";
WAIT FOR clk_period;
UR <= "111000101";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "111101110";
UI <= "010101000";
WAIT FOR clk_period;
UR <= "000010100";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "010100111";
WAIT FOR clk_period;
UR <= "001000111";
UI <= "010011000";
WAIT FOR clk_period;
UR <= "001010000";
UI <= "010000100";
WAIT FOR clk_period;
UR <= "001001110";
UI <= "001100011";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "000110001";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "111101001";
WAIT FOR clk_period;
UR <= "000000010";
UI <= "110111100";
WAIT FOR clk_period;
UR <= "111101000";
UI <= "110001111";
WAIT FOR clk_period;
UR <= "111010001";
UI <= "101100101";
WAIT FOR clk_period;
UR <= "110111101";
UI <= "101000000";
WAIT FOR clk_period;
UR <= "110101110";
UI <= "100100011";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "100010000";
WAIT FOR clk_period;
UR <= "110011110";
UI <= "100000001";
WAIT FOR clk_period;
UR <= "110011110";
UI <= "100000001";
WAIT FOR clk_period;
UR <= "110100100";
UI <= "100001100";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "100011101";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "100111101";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "101100100";
WAIT FOR clk_period;
UR <= "111101001";
UI <= "110010001";
WAIT FOR clk_period;
UR <= "000000011";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "000011011";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "001000100";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "001001101";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "001010000";
UI <= "010010010";
WAIT FOR clk_period;
UR <= "001000110";
UI <= "010100100";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "010101001";
WAIT FOR clk_period;
UR <= "000010100";
UI <= "010100111";
WAIT FOR clk_period;
UR <= "111101110";
UI <= "010011011";
WAIT FOR clk_period;
UR <= "111000100";
UI <= "010000110";
WAIT FOR clk_period;
UR <= "110011000";
UI <= "001101111";
WAIT FOR clk_period;
UR <= "101110010";
UI <= "001010111";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "000111111";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "000101111";
WAIT FOR clk_period;
UR <= "101000000";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "101010000";
UI <= "000100000";
WAIT FOR clk_period;
UR <= "101101100";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "110010010";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "111110000";
UI <= "001011101";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "001110101";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "010001011";
WAIT FOR clk_period;
UR <= "001001110";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "001001101";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "010110010";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010110000";
WAIT FOR clk_period;
UR <= "111101111";
UI <= "010100100";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "010010101";
WAIT FOR clk_period;
UR <= "110001010";
UI <= "010000001";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "001100111";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "001001011";
WAIT FOR clk_period;
UR <= "100110111";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "101000000";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "110001101";
UI <= "111101111";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "111100010";
WAIT FOR clk_period;
UR <= "000001001";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "001001010";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "010000010";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "010101101";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "011000100";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "011000100";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "010110010";
UI <= "111101000";
WAIT FOR clk_period;
UR <= "010001010";
UI <= "111110000";
WAIT FOR clk_period;
UR <= "001010100";
UI <= "111111001";
WAIT FOR clk_period;
UR <= "000010110";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "000001010";
WAIT FOR clk_period;
UR <= "110011000";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "101100100";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "100111010";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "100100011";
UI <= "000101111";
WAIT FOR clk_period;
UR <= "100010110";
UI <= "000110110";
WAIT FOR clk_period;
UR <= "100011010";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "100100110";
UI <= "000111111";
WAIT FOR clk_period;
UR <= "100111001";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101001110";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "101110010";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "101111010";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101111100";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "101111000";
UI <= "000011111";
WAIT FOR clk_period;
UR <= "101101110";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101100010";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "101001101";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "101001001";
UI <= "000011011";
WAIT FOR clk_period;
UR <= "101001101";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "101010111";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "101101010";
UI <= "001000010";
WAIT FOR clk_period;
UR <= "110000010";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "110011111";
UI <= "001100100";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "001110011";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "010000011";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "010001111";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010011011";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "010100011";
WAIT FOR clk_period;
UR <= "001001001";
UI <= "010100111";
WAIT FOR clk_period;
UR <= "001010111";
UI <= "010101011";
WAIT FOR clk_period;
UR <= "001100000";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "001100001";
UI <= "010101111";
WAIT FOR clk_period;
UR <= "001011111";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "001010110";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "001001000";
UI <= "010101011";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "010100111";
WAIT FOR clk_period;
UR <= "000011111";
UI <= "010100010";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "010011001";
WAIT FOR clk_period;
UR <= "111101011";
UI <= "010010000";
WAIT FOR clk_period;
UR <= "111001111";
UI <= "010000010";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "001110100";
WAIT FOR clk_period;
UR <= "110010111";
UI <= "001100101";
WAIT FOR clk_period;
UR <= "101111111";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "111101010";
WAIT FOR clk_period;
UR <= "101101110";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "111000100";
WAIT FOR clk_period;
UR <= "110010111";
UI <= "110101111";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "110011010";
WAIT FOR clk_period;
UR <= "111000101";
UI <= "110000100";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "101010110";
WAIT FOR clk_period;
UR <= "111111010";
UI <= "101000001";
WAIT FOR clk_period;
UR <= "000000001";
UI <= "100101101";
WAIT FOR clk_period;
UR <= "000000011";
UI <= "100011111";
WAIT FOR clk_period;
UR <= "111111110";
UI <= "100011000";
WAIT FOR clk_period;
UR <= "111110101";
UI <= "100011001";
WAIT FOR clk_period;
UR <= "111101000";
UI <= "100100010";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "100110111";
WAIT FOR clk_period;
UR <= "111001000";
UI <= "101010111";
WAIT FOR clk_period;
UR <= "110110101";
UI <= "101111100";
WAIT FOR clk_period;
UR <= "110100100";
UI <= "110101010";
WAIT FOR clk_period;
UR <= "110010100";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "110000111";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "101111101";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "101110011";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "101101100";
UI <= "001001110";
WAIT FOR clk_period;
UR <= "101101001";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000110111";
WAIT FOR clk_period;
UR <= "101101000";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "111101101";
WAIT FOR clk_period;
UR <= "101110100";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "110000000";
UI <= "110001101";
WAIT FOR clk_period;
UR <= "110001110";
UI <= "101100101";
WAIT FOR clk_period;
UR <= "110100000";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "110110110";
UI <= "100111100";
WAIT FOR clk_period;
UR <= "111001101";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "111100101";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "111111101";
UI <= "110000011";
WAIT FOR clk_period;
UR <= "000010010";
UI <= "110111011";
WAIT FOR clk_period;
UR <= "000100101";
UI <= "111111001";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "001101111";
WAIT FOR clk_period;
UR <= "000111101";
UI <= "010011101";
WAIT FOR clk_period;
UR <= "000111010";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "000110000";
UI <= "010111110";
WAIT FOR clk_period;
UR <= "000100000";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "000001101";
UI <= "010010010";
WAIT FOR clk_period;
UR <= "111111011";
UI <= "001100010";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "000101010";
WAIT FOR clk_period;
UR <= "111010110";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "111001100";
UI <= "110101111";
WAIT FOR clk_period;
UR <= "111000111";
UI <= "101111010";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "101010001";
WAIT FOR clk_period;
UR <= "111010110";
UI <= "100110110";
WAIT FOR clk_period;
UR <= "111100111";
UI <= "100101101";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "100110010";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "101000100";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "001011011";
UI <= "110000001";
WAIT FOR clk_period;
UR <= "001111001";
UI <= "110100110";
WAIT FOR clk_period;
UR <= "010010010";
UI <= "111001001";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "010110100";
UI <= "111111011";
WAIT FOR clk_period;
UR <= "010111110";
UI <= "000001001";
WAIT FOR clk_period;
UR <= "011000001";
UI <= "000001111";
WAIT FOR clk_period;
UR <= "010111111";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "010111010";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "010110001";
UI <= "111110111";
WAIT FOR clk_period;
UR <= "010101001";
UI <= "111101000";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "111010111";
WAIT FOR clk_period;
UR <= "010011011";
UI <= "111000111";
WAIT FOR clk_period;
UR <= "010010111";
UI <= "110111011";
WAIT FOR clk_period;
UR <= "010010101";
UI <= "110110001";
WAIT FOR clk_period;
UR <= "010010101";
UI <= "110101001";
WAIT FOR clk_period;
UR <= "010011000";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "010011100";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "010011110";
UI <= "110101101";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "110111010";
WAIT FOR clk_period;
UR <= "010100011";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "010100000";
UI <= "111111100";
WAIT FOR clk_period;
UR <= "010011001";
UI <= "000011001";
WAIT FOR clk_period;
UR <= "010010000";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "010000001";
UI <= "001011011";
WAIT FOR clk_period;
UR <= "001110001";
UI <= "001110110";
WAIT FOR clk_period;
UR <= "001011110";
UI <= "010001111";
WAIT FOR clk_period;
UR <= "001000110";
UI <= "010100010";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "111110111";
UI <= "010100100";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "010010100";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "001111111";
WAIT FOR clk_period;
UR <= "110100101";
UI <= "001100100";
WAIT FOR clk_period;
UR <= "110001101";
UI <= "001001001";
WAIT FOR clk_period;
UR <= "101111001";
UI <= "000110100";
WAIT FOR clk_period;
UR <= "101100111";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000011000";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101001011";
UI <= "000011000";
WAIT FOR clk_period;
UR <= "101001010";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "101001011";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101001110";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "001001101";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "001000111";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000111000";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101110110";
UI <= "111111111";
WAIT FOR clk_period;
UR <= "101111110";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "110000110";
UI <= "110110000";
WAIT FOR clk_period;
UR <= "110010011";
UI <= "110001011";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "101101010";
WAIT FOR clk_period;
UR <= "110110111";
UI <= "101010100";
WAIT FOR clk_period;
UR <= "111001110";
UI <= "101001000";
WAIT FOR clk_period;
UR <= "111101000";
UI <= "101000111";
WAIT FOR clk_period;
UR <= "000000101";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "000100100";
UI <= "101101011";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "110000111";
WAIT FOR clk_period;
UR <= "001011110";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "001111001";
UI <= "111000010";
WAIT FOR clk_period;
UR <= "010001100";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "010011100";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "010100100";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "010100100";
UI <= "111100101";
WAIT FOR clk_period;
UR <= "010011011";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "010001100";
UI <= "110111011";
WAIT FOR clk_period;
UR <= "001110110";
UI <= "110011110";
WAIT FOR clk_period;
UR <= "001011000";
UI <= "110000001";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "000010001";
UI <= "101010100";
WAIT FOR clk_period;
UR <= "111101001";
UI <= "101001011";
WAIT FOR clk_period;
UR <= "111000010";
UI <= "101001101";
WAIT FOR clk_period;
UR <= "110011100";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "101111001";
UI <= "101110011";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "110010011";
WAIT FOR clk_period;
UR <= "101001000";
UI <= "110110111";
WAIT FOR clk_period;
UR <= "100111011";
UI <= "111011111";
WAIT FOR clk_period;
UR <= "100111010";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "101000011";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "110011001";
UI <= "001001110";
WAIT FOR clk_period;
UR <= "111000111";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "111110101";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "000100111";
UI <= "000101011";
WAIT FOR clk_period;
UR <= "001010100";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "001111011";
UI <= "111111000";
WAIT FOR clk_period;
UR <= "010011010";
UI <= "111011101";
WAIT FOR clk_period;
UR <= "010101110";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "110101101";
WAIT FOR clk_period;
UR <= "010101110";
UI <= "110011000";
WAIT FOR clk_period;
UR <= "010011011";
UI <= "110000111";
WAIT FOR clk_period;
UR <= "001111101";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "001011001";
UI <= "101110000";
WAIT FOR clk_period;
UR <= "000101110";
UI <= "101101001";
WAIT FOR clk_period;
UR <= "000000011";
UI <= "101100101";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "101100011";
WAIT FOR clk_period;
UR <= "110110101";
UI <= "101101001";
WAIT FOR clk_period;
UR <= "110010100";
UI <= "101110001";
WAIT FOR clk_period;
UR <= "101111100";
UI <= "101111101";
WAIT FOR clk_period;
UR <= "101101100";
UI <= "110010001";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "110100110";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "111000010";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "101101000";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "101111001";
UI <= "001000111";
WAIT FOR clk_period;
UR <= "110000010";
UI <= "001100110";
WAIT FOR clk_period;
UR <= "110001110";
UI <= "010000010";
WAIT FOR clk_period;
UR <= "110011011";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "110101100";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "000011110";
UI <= "010011001";
WAIT FOR clk_period;
UR <= "001000100";
UI <= "010001001";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "001110011";
WAIT FOR clk_period;
UR <= "010010001";
UI <= "001011100";
WAIT FOR clk_period;
UR <= "010110010";
UI <= "001000101";
WAIT FOR clk_period;
UR <= "011001000";
UI <= "000101100";
WAIT FOR clk_period;
UR <= "011010100";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "011010011";
UI <= "111111110";
WAIT FOR clk_period;
UR <= "011000010";
UI <= "111101011";
WAIT FOR clk_period;
UR <= "010100100";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "001111011";
UI <= "111001010";
WAIT FOR clk_period;
UR <= "001001000";
UI <= "111000000";
WAIT FOR clk_period;
UR <= "000010001";
UI <= "110111010";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "110101000";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "101100010";
UI <= "111110001";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000111000";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "001100000";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "010001001";
WAIT FOR clk_period;
UR <= "110010101";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "110111010";
UI <= "011001001";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "011011001";
WAIT FOR clk_period;
UR <= "000000010";
UI <= "011011100";
WAIT FOR clk_period;
UR <= "000011111";
UI <= "011001111";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "010110011";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "010001001";
WAIT FOR clk_period;
UR <= "001000111";
UI <= "001010100";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "000011001";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "111011101";
WAIT FOR clk_period;
UR <= "000100001";
UI <= "110100100";
WAIT FOR clk_period;
UR <= "000001011";
UI <= "101110110";
WAIT FOR clk_period;
UR <= "111110011";
UI <= "101010110";
WAIT FOR clk_period;
UR <= "111011101";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "111001010";
UI <= "101001101";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "101100101";
WAIT FOR clk_period;
UR <= "110110101";
UI <= "110001100";
WAIT FOR clk_period;
UR <= "110110110";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "111111000";
WAIT FOR clk_period;
UR <= "111001100";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "111100011";
UI <= "001101000";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "010010011";
WAIT FOR clk_period;
UR <= "000011111";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "001000010";
UI <= "010111111";
WAIT FOR clk_period;
UR <= "001100101";
UI <= "010111011";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "010101000";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "010000111";
WAIT FOR clk_period;
UR <= "010111010";
UI <= "001011111";
WAIT FOR clk_period;
UR <= "011000111";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "011001000";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "010111100";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "111000001";
WAIT FOR clk_period;
UR <= "010000110";
UI <= "110101101";
WAIT FOR clk_period;
UR <= "001011011";
UI <= "110100100";
WAIT FOR clk_period;
UR <= "000101100";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "111111011";
UI <= "110110111";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "111001101";
WAIT FOR clk_period;
UR <= "110011110";
UI <= "111101000";
WAIT FOR clk_period;
UR <= "101111010";
UI <= "000000110";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "001011100";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "001110010";
WAIT FOR clk_period;
UR <= "101110111";
UI <= "010000000";
WAIT FOR clk_period;
UR <= "110010110";
UI <= "010001101";
WAIT FOR clk_period;
UR <= "110111001";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "000000101";
UI <= "010011011";
WAIT FOR clk_period;
UR <= "000100111";
UI <= "010011100";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "001011000";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "001100101";
UI <= "010010101";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "010010110";
WAIT FOR clk_period;
UR <= "001100110";
UI <= "010010100";
WAIT FOR clk_period;
UR <= "001011100";
UI <= "010010101";
WAIT FOR clk_period;
UR <= "001001101";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "010011101";
WAIT FOR clk_period;
UR <= "000101001";
UI <= "010100001";
WAIT FOR clk_period;
UR <= "000010111";
UI <= "010100111";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "111111101";
UI <= "010110100";
WAIT FOR clk_period;
UR <= "111110111";
UI <= "010111010";
WAIT FOR clk_period;
UR <= "111110111";
UI <= "010111100";
WAIT FOR clk_period;
UR <= "111111101";
UI <= "010111100";
WAIT FOR clk_period;
UR <= "000001001";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "001001100";
UI <= "010001011";
WAIT FOR clk_period;
UR <= "001101000";
UI <= "001110010";
WAIT FOR clk_period;
UR <= "010000001";
UI <= "001010111";
WAIT FOR clk_period;
UR <= "010011001";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "010101010";
UI <= "000011101";
WAIT FOR clk_period;
UR <= "010110011";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "010110100";
UI <= "111101001";
WAIT FOR clk_period;
UR <= "010101010";
UI <= "111010111";
WAIT FOR clk_period;
UR <= "010011000";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "001111010";
UI <= "111000101";
WAIT FOR clk_period;
UR <= "001010110";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "000101100";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "111011010";
WAIT FOR clk_period;
UR <= "111010001";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "110100100";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "101111101";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000101100";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "100110010";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "100101000";
UI <= "001011111";
WAIT FOR clk_period;
UR <= "100101000";
UI <= "001100101";
WAIT FOR clk_period;
UR <= "100101101";
UI <= "001100101";
WAIT FOR clk_period;
UR <= "100111000";
UI <= "001011111";
WAIT FOR clk_period;
UR <= "101000110";
UI <= "001010011";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "101100111";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "101111001";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "110000111";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "110010101";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "110100010";
UI <= "110101100";
WAIT FOR clk_period;
UR <= "110101101";
UI <= "110001111";
WAIT FOR clk_period;
UR <= "110111001";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "111000011";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "111001111";
UI <= "101011100";
WAIT FOR clk_period;
UR <= "111011101";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "111111110";
UI <= "101101011";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "101111011";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "110010000";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "001011111";
UI <= "110111001";
WAIT FOR clk_period;
UR <= "001111100";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "010011001";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "010110101";
UI <= "111100011";
WAIT FOR clk_period;
UR <= "011001110";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "011100011";
UI <= "111101000";
WAIT FOR clk_period;
UR <= "011110010";
UI <= "111100101";
WAIT FOR clk_period;
UR <= "011110101";
UI <= "111011110";
WAIT FOR clk_period;
UR <= "011110001";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "011100001";
UI <= "111010011";
WAIT FOR clk_period;
UR <= "011000110";
UI <= "111001111";
WAIT FOR clk_period;
UR <= "010100001";
UI <= "111001110";
WAIT FOR clk_period;
UR <= "001110011";
UI <= "111010011";
WAIT FOR clk_period;
UR <= "000111111";
UI <= "111011010";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "110100001";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "101111010";
UI <= "000010001";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "000101010";
WAIT FOR clk_period;
UR <= "101010111";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "101101100";
UI <= "000110111";
WAIT FOR clk_period;
UR <= "110001110";
UI <= "000111000";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "111110000";
UI <= "000101011";
WAIT FOR clk_period;
UR <= "000100110";
UI <= "000011011";
WAIT FOR clk_period;
UR <= "001011010";
UI <= "000001010";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "111110101";
WAIT FOR clk_period;
UR <= "010101010";
UI <= "111011101";
WAIT FOR clk_period;
UR <= "010111111";
UI <= "111000001";
WAIT FOR clk_period;
UR <= "011000110";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "010111101";
UI <= "110001011";
WAIT FOR clk_period;
UR <= "010100100";
UI <= "101110010";
WAIT FOR clk_period;
UR <= "010000000";
UI <= "101011110";
WAIT FOR clk_period;
UR <= "001010101";
UI <= "101001101";
WAIT FOR clk_period;
UR <= "000100100";
UI <= "101000111";
WAIT FOR clk_period;
UR <= "111110000";
UI <= "101001010";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "110010010";
UI <= "101101010";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "110000111";
WAIT FOR clk_period;
UR <= "101010010";
UI <= "110101010";
WAIT FOR clk_period;
UR <= "100111111";
UI <= "111001111";
WAIT FOR clk_period;
UR <= "100111000";
UI <= "111110101";
WAIT FOR clk_period;
UR <= "100111100";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "101000111";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "101110111";
UI <= "001000010";
WAIT FOR clk_period;
UR <= "110011000";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "000101010";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "000001110";
UI <= "111111000";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "111011110";
WAIT FOR clk_period;
UR <= "001011010";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "001111100";
UI <= "110111010";
WAIT FOR clk_period;
UR <= "010010111";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "010101011";
UI <= "111000010";
WAIT FOR clk_period;
UR <= "010111000";
UI <= "111011010";
WAIT FOR clk_period;
UR <= "010111011";
UI <= "111111100";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "010101000";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "001111101";
WAIT FOR clk_period;
UR <= "001110010";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "001001110";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "000100111";
UI <= "011000001";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "010111101";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "110110101";
UI <= "010010001";
WAIT FOR clk_period;
UR <= "110010110";
UI <= "001110000";
WAIT FOR clk_period;
UR <= "101111101";
UI <= "001001100";
WAIT FOR clk_period;
UR <= "101101100";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "101100010";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "101100100";
UI <= "000001110";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "000011100";
WAIT FOR clk_period;
UR <= "110000000";
UI <= "000110110";
WAIT FOR clk_period;
UR <= "110010100";
UI <= "001010111";
WAIT FOR clk_period;
UR <= "110101101";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "010011111";
WAIT FOR clk_period;
UR <= "111100101";
UI <= "010111000";
WAIT FOR clk_period;
UR <= "000000010";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "000011111";
UI <= "011000100";
WAIT FOR clk_period;
UR <= "000111101";
UI <= "010110100";
WAIT FOR clk_period;
UR <= "001011001";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "001110010";
UI <= "001101110";
WAIT FOR clk_period;
UR <= "010000110";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "010011001";
UI <= "000010001";
WAIT FOR clk_period;
UR <= "010100100";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "010101011";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "010101100";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "110110111";
WAIT FOR clk_period;
UR <= "010011100";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "010001101";
UI <= "111100011";
WAIT FOR clk_period;
UR <= "001111100";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "001011000";
UI <= "001101000";
WAIT FOR clk_period;
UR <= "001000110";
UI <= "010010001";
WAIT FOR clk_period;
UR <= "000111000";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "000101011";
UI <= "010111011";
WAIT FOR clk_period;
UR <= "000100001";
UI <= "010111000";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "010100100";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "001111111";
WAIT FOR clk_period;
UR <= "000001111";
UI <= "001001110";
WAIT FOR clk_period;
UR <= "000001100";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "000000101";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "111111100";
UI <= "110100010";
WAIT FOR clk_period;
UR <= "111101111";
UI <= "101110011";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "101001111";
WAIT FOR clk_period;
UR <= "111001110";
UI <= "100111010";
WAIT FOR clk_period;
UR <= "110110111";
UI <= "100110111";
WAIT FOR clk_period;
UR <= "110100000";
UI <= "101000101";
WAIT FOR clk_period;
UR <= "110001001";
UI <= "101100001";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "110000110";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "110110011";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "101011000";
UI <= "001000011";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "001101011";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "010001001";
WAIT FOR clk_period;
UR <= "110001100";
UI <= "010011101";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "010101001";
WAIT FOR clk_period;
UR <= "111000101";
UI <= "010101011";
WAIT FOR clk_period;
UR <= "111100101";
UI <= "010101010";
WAIT FOR clk_period;
UR <= "000000010";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "000100000";
UI <= "010010011";
WAIT FOR clk_period;
UR <= "000111001";
UI <= "010000110";
WAIT FOR clk_period;
UR <= "001010000";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "001100101";
UI <= "001101000";
WAIT FOR clk_period;
UR <= "001110100";
UI <= "001011010";
WAIT FOR clk_period;
UR <= "010000000";
UI <= "001001001";
WAIT FOR clk_period;
UR <= "010001011";
UI <= "000110110";
WAIT FOR clk_period;
UR <= "010010100";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "010011010";
UI <= "000001101";
WAIT FOR clk_period;
UR <= "010011111";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "111011000";
WAIT FOR clk_period;
UR <= "010100101";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "010100111";
UI <= "110100011";
WAIT FOR clk_period;
UR <= "010101000";
UI <= "110001111";
WAIT FOR clk_period;
UR <= "010101001";
UI <= "110000100";
WAIT FOR clk_period;
UR <= "010100111";
UI <= "110000000";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "110001000";
WAIT FOR clk_period;
UR <= "010100011";
UI <= "110011100";
WAIT FOR clk_period;
UR <= "010011111";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "010011001";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "010010001";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "001111101";
UI <= "001111011";
WAIT FOR clk_period;
UR <= "001110001";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "001100010";
UI <= "011000010";
WAIT FOR clk_period;
UR <= "001010001";
UI <= "011010001";
WAIT FOR clk_period;
UR <= "000111101";
UI <= "011001100";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "010110011";
WAIT FOR clk_period;
UR <= "000010101";
UI <= "010001100";
WAIT FOR clk_period;
UR <= "000000000";
UI <= "001010101";
WAIT FOR clk_period;
UR <= "111101110";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "111011101";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "110011001";
WAIT FOR clk_period;
UR <= "111001010";
UI <= "101101001";
WAIT FOR clk_period;
UR <= "111001000";
UI <= "101001001";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "100111101";
WAIT FOR clk_period;
UR <= "111010110";
UI <= "101001000";
WAIT FOR clk_period;
UR <= "111100010";
UI <= "101101000";
WAIT FOR clk_period;
UR <= "111110001";
UI <= "110011001";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "000010101";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "000100100";
UI <= "001010111";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "010001011";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "011000011";
WAIT FOR clk_period;
UR <= "000101100";
UI <= "010111111";
WAIT FOR clk_period;
UR <= "000100000";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "000010001";
UI <= "001111001";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "111011101";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "110000100";
WAIT FOR clk_period;
UR <= "111001101";
UI <= "101010111";
WAIT FOR clk_period;
UR <= "111010000";
UI <= "100110111";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "100101010";
WAIT FOR clk_period;
UR <= "111101011";
UI <= "100101111";
WAIT FOR clk_period;
UR <= "000000001";
UI <= "101000010";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "000111110";
UI <= "110000110";
WAIT FOR clk_period;
UR <= "001011111";
UI <= "110101100";
WAIT FOR clk_period;
UR <= "001111111";
UI <= "111010000";
WAIT FOR clk_period;
UR <= "010011100";
UI <= "111101010";
WAIT FOR clk_period;
UR <= "010110100";
UI <= "111111011";
WAIT FOR clk_period;
UR <= "011000111";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "011010001";
UI <= "111111101";
WAIT FOR clk_period;
UR <= "011010111";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "011010110";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "011001110";
UI <= "111010001";
WAIT FOR clk_period;
UR <= "011000011";
UI <= "111000101";
WAIT FOR clk_period;
UR <= "010110001";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "010100000";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "010001011";
UI <= "111000111";
WAIT FOR clk_period;
UR <= "001110110";
UI <= "111011010";
WAIT FOR clk_period;
UR <= "001100101";
UI <= "111110101";
WAIT FOR clk_period;
UR <= "001010100";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "001000110";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "001011111";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "010000010";
WAIT FOR clk_period;
UR <= "000110000";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "000110000";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "000110001";
UI <= "011001111";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "011010000";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "011001101";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "000110011";
UI <= "010111011";
WAIT FOR clk_period;
UR <= "000110001";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "010011111";
WAIT FOR clk_period;
UR <= "000100000";
UI <= "010010010";
WAIT FOR clk_period;
UR <= "000010100";
UI <= "010000011";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "001110101";
WAIT FOR clk_period;
UR <= "111101110";
UI <= "001100111";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "001011001";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "001001011";
WAIT FOR clk_period;
UR <= "110100101";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "110000111";
UI <= "000110111";
WAIT FOR clk_period;
UR <= "101101011";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "100110110";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "100100001";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "100010011";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "100001100";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "100001111";
UI <= "000101000";
WAIT FOR clk_period;
UR <= "100011110";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "100110110";
UI <= "000110000";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000110000";
WAIT FOR clk_period;
UR <= "110000110";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "110111010";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "111101111";
UI <= "000011111";
WAIT FOR clk_period;
UR <= "000100101";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "001010111";
UI <= "000000101";
WAIT FOR clk_period;
UR <= "010000001";
UI <= "111110101";
WAIT FOR clk_period;
UR <= "010100001";
UI <= "111100101";
WAIT FOR clk_period;
UR <= "010110010";
UI <= "111010100";
WAIT FOR clk_period;
UR <= "010110100";
UI <= "111000100";
WAIT FOR clk_period;
UR <= "010101000";
UI <= "110110111";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "110101001";
WAIT FOR clk_period;
UR <= "001101101";
UI <= "110100000";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "110010101";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "110001100";
WAIT FOR clk_period;
UR <= "111110100";
UI <= "110000011";
WAIT FOR clk_period;
UR <= "111010110";
UI <= "101110111";
WAIT FOR clk_period;
UR <= "110111110";
UI <= "101101100";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "101010001";
WAIT FOR clk_period;
UR <= "110111011";
UI <= "101000101";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "100111101";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "100110110";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "100110100";
WAIT FOR clk_period;
UR <= "111110101";
UI <= "100111001";
WAIT FOR clk_period;
UR <= "111110111";
UI <= "101000100";
WAIT FOR clk_period;
UR <= "111101111";
UI <= "101011001";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "101110001";
WAIT FOR clk_period;
UR <= "110111110";
UI <= "110010000";
WAIT FOR clk_period;
UR <= "110011100";
UI <= "110110001";
WAIT FOR clk_period;
UR <= "101111001";
UI <= "111010011";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "101000011";
UI <= "000001110";
WAIT FOR clk_period;
UR <= "100110111";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "100111100";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000111000";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "110100101";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "000010110";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "001001110";
UI <= "111110111";
WAIT FOR clk_period;
UR <= "001111111";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "010100011";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "010110101";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "010110111";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "111001010";
WAIT FOR clk_period;
UR <= "010000110";
UI <= "111010010";
WAIT FOR clk_period;
UR <= "001011000";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "000100011";
UI <= "111110011";
WAIT FOR clk_period;
UR <= "111100111";
UI <= "000000100";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101111000";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101001011";
UI <= "000110110";
WAIT FOR clk_period;
UR <= "100100111";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "100001111";
UI <= "001000111";
WAIT FOR clk_period;
UR <= "100000001";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "011111111";
UI <= "001000101";
WAIT FOR clk_period;
UR <= "100001000";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "100011001";
UI <= "000111000";
WAIT FOR clk_period;
UR <= "100110011";
UI <= "000101111";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "110011101";
UI <= "000011001";
WAIT FOR clk_period;
UR <= "111000110";
UI <= "000010010";
WAIT FOR clk_period;
UR <= "111110001";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "000000100";
WAIT FOR clk_period;
UR <= "001000100";
UI <= "111111100";
WAIT FOR clk_period;
UR <= "001101000";
UI <= "111110100";
WAIT FOR clk_period;
UR <= "010001010";
UI <= "111101001";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "111011111";
WAIT FOR clk_period;
UR <= "010110101";
UI <= "111010001";
WAIT FOR clk_period;
UR <= "011000000";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "011000011";
UI <= "110111011";
WAIT FOR clk_period;
UR <= "011000001";
UI <= "110110100";
WAIT FOR clk_period;
UR <= "010111000";
UI <= "110101111";
WAIT FOR clk_period;
UR <= "010101110";
UI <= "110110000";
WAIT FOR clk_period;
UR <= "010100010";
UI <= "110110110";
WAIT FOR clk_period;
UR <= "010010101";
UI <= "111000000";
WAIT FOR clk_period;
UR <= "010001101";
UI <= "111010001";
WAIT FOR clk_period;
UR <= "010001001";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "010000110";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "010001010";
UI <= "000111100";
WAIT FOR clk_period;
UR <= "010000111";
UI <= "001011011";
WAIT FOR clk_period;
UR <= "010000001";
UI <= "001110101";
WAIT FOR clk_period;
UR <= "001110010";
UI <= "010001100";
WAIT FOR clk_period;
UR <= "001011011";
UI <= "010011111";
WAIT FOR clk_period;
UR <= "000111001";
UI <= "010101001";
WAIT FOR clk_period;
UR <= "000001110";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "111011110";
UI <= "010101001";
WAIT FOR clk_period;
UR <= "110101010";
UI <= "010011101";
WAIT FOR clk_period;
UR <= "101111101";
UI <= "010001100";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "001111000";
WAIT FOR clk_period;
UR <= "100110111";
UI <= "001100000";
WAIT FOR clk_period;
UR <= "100101101";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "100110101";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "101010010";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "110111011";
UI <= "111110000";
WAIT FOR clk_period;
UR <= "111111100";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "001000000";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "001111011";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "010101010";
UI <= "111010101";
WAIT FOR clk_period;
UR <= "011000011";
UI <= "111010111";
WAIT FOR clk_period;
UR <= "011001001";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "010110101";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "010001110";
UI <= "111101001";
WAIT FOR clk_period;
UR <= "001010101";
UI <= "111110010";
WAIT FOR clk_period;
UR <= "000010010";
UI <= "111111010";
WAIT FOR clk_period;
UR <= "111001101";
UI <= "000000100";
WAIT FOR clk_period;
UR <= "110001110";
UI <= "000001101";
WAIT FOR clk_period;
UR <= "101011100";
UI <= "000011000";
WAIT FOR clk_period;
UR <= "100111101";
UI <= "000011110";
WAIT FOR clk_period;
UR <= "100110110";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101000110";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "101101011";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "111100011";
UI <= "000101100";
WAIT FOR clk_period;
UR <= "000101000";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "001101000";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "010011101";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "011000010";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "011010010";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "011001101";
UI <= "110101011";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "110001100";
WAIT FOR clk_period;
UR <= "010001101";
UI <= "101101110";
WAIT FOR clk_period;
UR <= "001011101";
UI <= "101010111";
WAIT FOR clk_period;
UR <= "000101000";
UI <= "101000111";
WAIT FOR clk_period;
UR <= "111110111";
UI <= "101000000";
WAIT FOR clk_period;
UR <= "111001101";
UI <= "101000110";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "101010100";
WAIT FOR clk_period;
UR <= "110100001";
UI <= "101101111";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "110010011";
WAIT FOR clk_period;
UR <= "110110000";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "111101111";
WAIT FOR clk_period;
UR <= "111101001";
UI <= "000100000";
WAIT FOR clk_period;
UR <= "000001010";
UI <= "001001110";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "001111001";
WAIT FOR clk_period;
UR <= "001000010";
UI <= "010011100";
WAIT FOR clk_period;
UR <= "001010001";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "001010111";
UI <= "011000100";
WAIT FOR clk_period;
UR <= "001010010";
UI <= "011001010";
WAIT FOR clk_period;
UR <= "001001000";
UI <= "011001000";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "011000001";
WAIT FOR clk_period;
UR <= "000100111";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "000011001";
UI <= "010101010";
WAIT FOR clk_period;
UR <= "000010000";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "000001101";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "010010000";
WAIT FOR clk_period;
UR <= "000011110";
UI <= "010010010";
WAIT FOR clk_period;
UR <= "000101111";
UI <= "010010110";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "001010001";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "001011101";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "001011110";
UI <= "010110011";
WAIT FOR clk_period;
UR <= "001011000";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "001000101";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "000101000";
UI <= "010100100";
WAIT FOR clk_period;
UR <= "000000011";
UI <= "010010011";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "001111110";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "001101000";
WAIT FOR clk_period;
UR <= "110000111";
UI <= "001010010";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101001000";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "101001100";
UI <= "000100000";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "101111100";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "110100000";
UI <= "001000010";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "001010111";
WAIT FOR clk_period;
UR <= "111110001";
UI <= "001101110";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "010000101";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "010011001";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "010101000";
WAIT FOR clk_period;
UR <= "000111110";
UI <= "010110000";
WAIT FOR clk_period;
UR <= "000110001";
UI <= "010110010";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "010011111";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "010001100";
WAIT FOR clk_period;
UR <= "110101011";
UI <= "001110101";
WAIT FOR clk_period;
UR <= "110000101";
UI <= "001011011";
WAIT FOR clk_period;
UR <= "101100111";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "101000011";
UI <= "000000110";
WAIT FOR clk_period;
UR <= "101000011";
UI <= "111101111";
WAIT FOR clk_period;
UR <= "101001110";
UI <= "111011000";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "111000001";
WAIT FOR clk_period;
UR <= "101111010";
UI <= "110110000";
WAIT FOR clk_period;
UR <= "110011001";
UI <= "110011110";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "110001101";
WAIT FOR clk_period;
UR <= "111010100";
UI <= "101111010";
WAIT FOR clk_period;
UR <= "111101010";
UI <= "101101001";
WAIT FOR clk_period;
UR <= "111111011";
UI <= "101010111";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "101000111";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "100111010";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "100110000";
WAIT FOR clk_period;
UR <= "111110110";
UI <= "100101100";
WAIT FOR clk_period;
UR <= "111101000";
UI <= "100101100";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "100110110";
WAIT FOR clk_period;
UR <= "111001000";
UI <= "101000110";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "101011110";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "101111100";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "110011110";
WAIT FOR clk_period;
UR <= "110011111";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "110011001";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "110010010";
UI <= "000000111";
WAIT FOR clk_period;
UR <= "110001010";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101111110";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101110011";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "100110110";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "100101011";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "100101000";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "100101110";
UI <= "000001010";
WAIT FOR clk_period;
UR <= "100111010";
UI <= "000010000";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000011101";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "110010011";
UI <= "001001110";
WAIT FOR clk_period;
UR <= "110111011";
UI <= "001101110";
WAIT FOR clk_period;
UR <= "111100001";
UI <= "010001100";
WAIT FOR clk_period;
UR <= "000000101";
UI <= "010100100";
WAIT FOR clk_period;
UR <= "000100001";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "010111111";
WAIT FOR clk_period;
UR <= "000111110";
UI <= "010111000";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "000110000";
UI <= "010000110";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "001011011";
WAIT FOR clk_period;
UR <= "000000100";
UI <= "000101010";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "111110111";
WAIT FOR clk_period;
UR <= "111010110";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "111000110";
UI <= "110010100";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "101101111";
WAIT FOR clk_period;
UR <= "111000010";
UI <= "101010100";
WAIT FOR clk_period;
UR <= "111010000";
UI <= "101000110";
WAIT FOR clk_period;
UR <= "111101000";
UI <= "101000101";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "101010000";
WAIT FOR clk_period;
UR <= "000101011";
UI <= "101100100";
WAIT FOR clk_period;
UR <= "001010011";
UI <= "101111110";
WAIT FOR clk_period;
UR <= "001110101";
UI <= "110011011";
WAIT FOR clk_period;
UR <= "010010010";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "111010000";
WAIT FOR clk_period;
UR <= "010110000";
UI <= "111100010";
WAIT FOR clk_period;
UR <= "010101100";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "010100000";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "001101010";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "001000111";
UI <= "110111110";
WAIT FOR clk_period;
UR <= "000100001";
UI <= "110100011";
WAIT FOR clk_period;
UR <= "111111110";
UI <= "110000110";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "111000010";
UI <= "101001100";
WAIT FOR clk_period;
UR <= "110101101";
UI <= "100110011";
WAIT FOR clk_period;
UR <= "110100000";
UI <= "100100011";
WAIT FOR clk_period;
UR <= "110011000";
UI <= "100011001";
WAIT FOR clk_period;
UR <= "110011001";
UI <= "100010101";
WAIT FOR clk_period;
UR <= "110100001";
UI <= "100011011";
WAIT FOR clk_period;
UR <= "110101110";
UI <= "100101000";
WAIT FOR clk_period;
UR <= "110111110";
UI <= "100111101";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "101011011";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "101111101";
WAIT FOR clk_period;
UR <= "111111100";
UI <= "110101001";
WAIT FOR clk_period;
UR <= "000010000";
UI <= "111010100";
WAIT FOR clk_period;
UR <= "000100010";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "000110000";
UI <= "000101011";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "001010100";
WAIT FOR clk_period;
UR <= "000111110";
UI <= "001110110";
WAIT FOR clk_period;
UR <= "000111011";
UI <= "010010010";
WAIT FOR clk_period;
UR <= "000110000";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "000011110";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "111101010";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "111001000";
UI <= "010010100";
WAIT FOR clk_period;
UR <= "110101000";
UI <= "001111110";
WAIT FOR clk_period;
UR <= "110001000";
UI <= "001100011";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101001100";
UI <= "000011101";
WAIT FOR clk_period;
UR <= "101000110";
UI <= "000001101";
WAIT FOR clk_period;
UR <= "101000111";
UI <= "000000100";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101110110";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "101110110";
UI <= "000110000";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "101001111";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "100111110";
UI <= "001001001";
WAIT FOR clk_period;
UR <= "100101110";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "100100100";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "100100100";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "100101111";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101001001";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "110100000";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "000000001";
WAIT FOR clk_period;
UR <= "000010011";
UI <= "111110111";
WAIT FOR clk_period;
UR <= "001001100";
UI <= "111101111";
WAIT FOR clk_period;
UR <= "001111100";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "010100001";
UI <= "111100010";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "111011100";
WAIT FOR clk_period;
UR <= "010111001";
UI <= "111011010";
WAIT FOR clk_period;
UR <= "010101010";
UI <= "111011010";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "111011100";
WAIT FOR clk_period;
UR <= "001011100";
UI <= "111100001";
WAIT FOR clk_period;
UR <= "000100110";
UI <= "111101011";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "111110101";
WAIT FOR clk_period;
UR <= "110110010";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "101111110";
UI <= "000010010";
WAIT FOR clk_period;
UR <= "101010010";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "100110011";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "100100010";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "100011010";
UI <= "001010000";
WAIT FOR clk_period;
UR <= "100100000";
UI <= "001011000";
WAIT FOR clk_period;
UR <= "100101011";
UI <= "001011010";
WAIT FOR clk_period;
UR <= "100111011";
UI <= "001011001";
WAIT FOR clk_period;
UR <= "101001101";
UI <= "001001110";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "000111111";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "101111101";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "110000111";
UI <= "111111010";
WAIT FOR clk_period;
UR <= "110001110";
UI <= "111011101";
WAIT FOR clk_period;
UR <= "110010101";
UI <= "111000000";
WAIT FOR clk_period;
UR <= "110011100";
UI <= "110100110";
WAIT FOR clk_period;
UR <= "110100110";
UI <= "110001101";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "101101000";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "101011101";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "101011010";
WAIT FOR clk_period;
UR <= "000000110";
UI <= "101011001";
WAIT FOR clk_period;
UR <= "000100010";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "000111101";
UI <= "101101010";
WAIT FOR clk_period;
UR <= "001011010";
UI <= "101111010";
WAIT FOR clk_period;
UR <= "001110001";
UI <= "110001111";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "110101000";
WAIT FOR clk_period;
UR <= "010011010";
UI <= "111000100";
WAIT FOR clk_period;
UR <= "010100110";
UI <= "111100011";
WAIT FOR clk_period;
UR <= "010101111";
UI <= "000000101";
WAIT FOR clk_period;
UR <= "010110010";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "010101110";
UI <= "001001001";
WAIT FOR clk_period;
UR <= "010100100";
UI <= "001101000";
WAIT FOR clk_period;
UR <= "010010100";
UI <= "010000100";
WAIT FOR clk_period;
UR <= "001111100";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "001011101";
UI <= "010101000";
WAIT FOR clk_period;
UR <= "000111000";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "000001110";
UI <= "010101010";
WAIT FOR clk_period;
UR <= "111011111";
UI <= "010100001";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "010001111";
WAIT FOR clk_period;
UR <= "110001010";
UI <= "001111001";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "001011111";
WAIT FOR clk_period;
UR <= "101001100";
UI <= "001000111";
WAIT FOR clk_period;
UR <= "100111111";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101000001";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101010011";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101110011";
UI <= "000001111";
WAIT FOR clk_period;
UR <= "110100000";
UI <= "000001110";
WAIT FOR clk_period;
UR <= "111010100";
UI <= "000010001";
WAIT FOR clk_period;
UR <= "000001101";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "001000100";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "001110110";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "010011101";
UI <= "000001010";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "111111000";
WAIT FOR clk_period;
UR <= "010111101";
UI <= "111011110";
WAIT FOR clk_period;
UR <= "010110011";
UI <= "110111100";
WAIT FOR clk_period;
UR <= "010011100";
UI <= "110010101";
WAIT FOR clk_period;
UR <= "001110110";
UI <= "101101111";
WAIT FOR clk_period;
UR <= "001001011";
UI <= "101001101";
WAIT FOR clk_period;
UR <= "000011100";
UI <= "100110010";
WAIT FOR clk_period;
UR <= "111110011";
UI <= "100100101";
WAIT FOR clk_period;
UR <= "111001111";
UI <= "100101000";
WAIT FOR clk_period;
UR <= "110110110";
UI <= "100111110";
WAIT FOR clk_period;
UR <= "110101110";
UI <= "101100011";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "110010111";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "111010110";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "111111000";
UI <= "001010110";
WAIT FOR clk_period;
UR <= "000010110";
UI <= "010001101";
WAIT FOR clk_period;
UR <= "000110001";
UI <= "010110010";
WAIT FOR clk_period;
UR <= "001000101";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "001001100";
UI <= "011000011";
WAIT FOR clk_period;
UR <= "001000111";
UI <= "010101000";
WAIT FOR clk_period;
UR <= "000111010";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "000100011";
UI <= "001000010";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "111010001";
UI <= "110000011";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "101010111";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "100111110";
WAIT FOR clk_period;
UR <= "110111010";
UI <= "100111100";
WAIT FOR clk_period;
UR <= "111000101";
UI <= "101001111";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "101110110";
WAIT FOR clk_period;
UR <= "111111000";
UI <= "110101101";
WAIT FOR clk_period;
UR <= "000010100";
UI <= "111101100";
WAIT FOR clk_period;
UR <= "000101110";
UI <= "000101101";
WAIT FOR clk_period;
UR <= "001000010";
UI <= "001101100";
WAIT FOR clk_period;
UR <= "001001010";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "001001000";
UI <= "011000000";
WAIT FOR clk_period;
UR <= "000111001";
UI <= "011010011";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "011010011";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "011000001";
WAIT FOR clk_period;
UR <= "111010000";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "110100100";
UI <= "010000000";
WAIT FOR clk_period;
UR <= "101111110";
UI <= "001011001";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000110111";
WAIT FOR clk_period;
UR <= "101001100";
UI <= "000011100";
WAIT FOR clk_period;
UR <= "101000110";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "101001110";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "000010000";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "111010001";
UI <= "001011100";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "001111100";
WAIT FOR clk_period;
UR <= "000011010";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "000110110";
UI <= "010110000";
WAIT FOR clk_period;
UR <= "001001010";
UI <= "010111111";
WAIT FOR clk_period;
UR <= "001010011";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "001010011";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "001001100";
UI <= "011000000";
WAIT FOR clk_period;
UR <= "001000001";
UI <= "010110110";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "010101010";
WAIT FOR clk_period;
UR <= "000101001";
UI <= "010100001";
WAIT FOR clk_period;
UR <= "000100000";
UI <= "010010111";
WAIT FOR clk_period;
UR <= "000011011";
UI <= "010010010";
WAIT FOR clk_period;
UR <= "000011011";
UI <= "010010011";
WAIT FOR clk_period;
UR <= "000100001";
UI <= "010010100";
WAIT FOR clk_period;
UR <= "000101001";
UI <= "010011010";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "010100000";
WAIT FOR clk_period;
UR <= "000111110";
UI <= "010100111";
WAIT FOR clk_period;
UR <= "001000011";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "001000110";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "001000010";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "000110110";
UI <= "010100111";
WAIT FOR clk_period;
UR <= "000100100";
UI <= "010011111";
WAIT FOR clk_period;
UR <= "000001011";
UI <= "010010000";
WAIT FOR clk_period;
UR <= "111101110";
UI <= "010000000";
WAIT FOR clk_period;
UR <= "111001101";
UI <= "001101111";
WAIT FOR clk_period;
UR <= "110101101";
UI <= "001011110";
WAIT FOR clk_period;
UR <= "110001110";
UI <= "001001100";
WAIT FOR clk_period;
UR <= "101110011";
UI <= "000111100";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101001101";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "101000100";
UI <= "000011010";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "000010101";
WAIT FOR clk_period;
UR <= "101000010";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "101001001";
UI <= "000010100";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "000011001";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "000011111";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000101110";
WAIT FOR clk_period;
UR <= "101101000";
UI <= "000110101";
WAIT FOR clk_period;
UR <= "101101001";
UI <= "000111100";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "001000100";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "101010111";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "101101011";
UI <= "000000100";
WAIT FOR clk_period;
UR <= "101111001";
UI <= "111110000";
WAIT FOR clk_period;
UR <= "110001001";
UI <= "111011000";
WAIT FOR clk_period;
UR <= "110011101";
UI <= "111000000";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "110100111";
WAIT FOR clk_period;
UR <= "111000010";
UI <= "110001110";
WAIT FOR clk_period;
UR <= "111010011";
UI <= "101110100";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "101011011";
WAIT FOR clk_period;
UR <= "111101100";
UI <= "101000111";
WAIT FOR clk_period;
UR <= "111110001";
UI <= "100110100";
WAIT FOR clk_period;
UR <= "111110100";
UI <= "100100110";
WAIT FOR clk_period;
UR <= "111110100";
UI <= "100011111";
WAIT FOR clk_period;
UR <= "111101110";
UI <= "100011110";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "100100101";
WAIT FOR clk_period;
UR <= "111011011";
UI <= "100110110";
WAIT FOR clk_period;
UR <= "111001111";
UI <= "101001110";
WAIT FOR clk_period;
UR <= "111000011";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "110110111";
UI <= "110010001";
WAIT FOR clk_period;
UR <= "110101001";
UI <= "110111001";
WAIT FOR clk_period;
UR <= "110011101";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "110010000";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "110000101";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101111010";
UI <= "000110011";
WAIT FOR clk_period;
UR <= "101110000";
UI <= "000111110";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000111010";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "000101011";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000010001";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "111110001";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "101101110";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "110000011";
WAIT FOR clk_period;
UR <= "110011000";
UI <= "101100111";
WAIT FOR clk_period;
UR <= "110110111";
UI <= "101010100";
WAIT FOR clk_period;
UR <= "111011001";
UI <= "101001100";
WAIT FOR clk_period;
UR <= "000000010";
UI <= "101010000";
WAIT FOR clk_period;
UR <= "000101010";
UI <= "101011110";
WAIT FOR clk_period;
UR <= "001010001";
UI <= "101110100";
WAIT FOR clk_period;
UR <= "001110100";
UI <= "110001111";
WAIT FOR clk_period;
UR <= "010010001";
UI <= "110101010";
WAIT FOR clk_period;
UR <= "010100101";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "010101111";
UI <= "111011000";
WAIT FOR clk_period;
UR <= "010101110";
UI <= "111100100";
WAIT FOR clk_period;
UR <= "010100001";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "010001100";
UI <= "111011111";
WAIT FOR clk_period;
UR <= "001101110";
UI <= "111010000";
WAIT FOR clk_period;
UR <= "001001010";
UI <= "110111010";
WAIT FOR clk_period;
UR <= "000100111";
UI <= "110100000";
WAIT FOR clk_period;
UR <= "000000110";
UI <= "110000111";
WAIT FOR clk_period;
UR <= "111101010";
UI <= "101101111";
WAIT FOR clk_period;
UR <= "111010100";
UI <= "101011110";
WAIT FOR clk_period;
UR <= "111001010";
UI <= "101010001";
WAIT FOR clk_period;
UR <= "111001011";
UI <= "101001111";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "101010011";
WAIT FOR clk_period;
UR <= "111101011";
UI <= "101011111";
WAIT FOR clk_period;
UR <= "000001001";
UI <= "101110011";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "110001000";
WAIT FOR clk_period;
UR <= "001010010";
UI <= "110100000";
WAIT FOR clk_period;
UR <= "001110111";
UI <= "110111000";
WAIT FOR clk_period;
UR <= "010011010";
UI <= "111001110";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "111100010";
WAIT FOR clk_period;
UR <= "011001100";
UI <= "111110010";
WAIT FOR clk_period;
UR <= "011010111";
UI <= "111111101";
WAIT FOR clk_period;
UR <= "011011110";
UI <= "000000011";
WAIT FOR clk_period;
UR <= "011011100";
UI <= "000000100";
WAIT FOR clk_period;
UR <= "011010010";
UI <= "000000010";
WAIT FOR clk_period;
UR <= "011000100";
UI <= "111111001";
WAIT FOR clk_period;
UR <= "010110011";
UI <= "111101101";
WAIT FOR clk_period;
UR <= "010011110";
UI <= "111011101";
WAIT FOR clk_period;
UR <= "010001001";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "001110011";
UI <= "110110011";
WAIT FOR clk_period;
UR <= "001011100";
UI <= "110011010";
WAIT FOR clk_period;
UR <= "001000111";
UI <= "110000100";
WAIT FOR clk_period;
UR <= "000110001";
UI <= "101101111";
WAIT FOR clk_period;
UR <= "000011101";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "000000111";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "111110010";
UI <= "101010001";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "101010101";
WAIT FOR clk_period;
UR <= "111000110";
UI <= "101100010";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "101111000";
WAIT FOR clk_period;
UR <= "110011100";
UI <= "110010101";
WAIT FOR clk_period;
UR <= "110001001";
UI <= "110110101";
WAIT FOR clk_period;
UR <= "101111001";
UI <= "111011001";
WAIT FOR clk_period;
UR <= "101101101";
UI <= "111111011";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "000011001";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "001000011";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "001001011";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "001000011";
WAIT FOR clk_period;
UR <= "101011111";
UI <= "000110110";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101100011";
UI <= "000011101";
WAIT FOR clk_period;
UR <= "101100010";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "101100001";
UI <= "000010011";
WAIT FOR clk_period;
UR <= "101100000";
UI <= "000011001";
WAIT FOR clk_period;
UR <= "101011101";
UI <= "000100011";
WAIT FOR clk_period;
UR <= "101011001";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101010111";
UI <= "001000011";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "001010011";
WAIT FOR clk_period;
UR <= "101010101";
UI <= "001011111";
WAIT FOR clk_period;
UR <= "101010110";
UI <= "001100010";
WAIT FOR clk_period;
UR <= "101011010";
UI <= "001011010";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "101100101";
UI <= "000101001";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "000000000";
WAIT FOR clk_period;
UR <= "101111011";
UI <= "111010010";
WAIT FOR clk_period;
UR <= "110000111";
UI <= "110100100";
WAIT FOR clk_period;
UR <= "110010110";
UI <= "101111001";
WAIT FOR clk_period;
UR <= "110100110";
UI <= "101010111";
WAIT FOR clk_period;
UR <= "110110110";
UI <= "101000011";
WAIT FOR clk_period;
UR <= "111001000";
UI <= "100111111";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "101001011";
WAIT FOR clk_period;
UR <= "111101010";
UI <= "101101010";
WAIT FOR clk_period;
UR <= "111111001";
UI <= "110010110";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "000010101";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "000011110";
UI <= "001000001";
WAIT FOR clk_period;
UR <= "000100110";
UI <= "001110100";
WAIT FOR clk_period;
UR <= "000101011";
UI <= "010011100";
WAIT FOR clk_period;
UR <= "000101100";
UI <= "010110100";
WAIT FOR clk_period;
UR <= "000101001";
UI <= "010111000";
WAIT FOR clk_period;
UR <= "000100110";
UI <= "010101011";
WAIT FOR clk_period;
UR <= "000011111";
UI <= "010001110";
WAIT FOR clk_period;
UR <= "000010101";
UI <= "001100001";
WAIT FOR clk_period;
UR <= "000001010";
UI <= "000101100";
WAIT FOR clk_period;
UR <= "111111111";
UI <= "111110000";
WAIT FOR clk_period;
UR <= "111110001";
UI <= "110110101";
WAIT FOR clk_period;
UR <= "111100110";
UI <= "101111110";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "101010000";
WAIT FOR clk_period;
UR <= "111001100";
UI <= "100101011";
WAIT FOR clk_period;
UR <= "111000001";
UI <= "100010011";
WAIT FOR clk_period;
UR <= "110111010";
UI <= "100001010";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "100001100";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "100010110";
WAIT FOR clk_period;
UR <= "110110011";
UI <= "100101000";
WAIT FOR clk_period;
UR <= "110111001";
UI <= "101000000";
WAIT FOR clk_period;
UR <= "111000100";
UI <= "101011001";
WAIT FOR clk_period;
UR <= "111010100";
UI <= "101110101";
WAIT FOR clk_period;
UR <= "111101001";
UI <= "110001100";
WAIT FOR clk_period;
UR <= "000000001";
UI <= "110011111";
WAIT FOR clk_period;
UR <= "000011110";
UI <= "110110001";
WAIT FOR clk_period;
UR <= "000111100";
UI <= "110111101";
WAIT FOR clk_period;
UR <= "001011001";
UI <= "111000101";
WAIT FOR clk_period;
UR <= "001110110";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "111001101";
WAIT FOR clk_period;
UR <= "010100011";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "010110011";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "010111100";
UI <= "111001000";
WAIT FOR clk_period;
UR <= "010111111";
UI <= "111000110";
WAIT FOR clk_period;
UR <= "010111110";
UI <= "111000100";
WAIT FOR clk_period;
UR <= "010111001";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "010110000";
UI <= "111000100";
WAIT FOR clk_period;
UR <= "010100101";
UI <= "111000111";
WAIT FOR clk_period;
UR <= "010011110";
UI <= "111001110";
WAIT FOR clk_period;
UR <= "010010101";
UI <= "111011000";
WAIT FOR clk_period;
UR <= "010001111";
UI <= "111100101";
WAIT FOR clk_period;
UR <= "010001001";
UI <= "111110111";
WAIT FOR clk_period;
UR <= "010000110";
UI <= "000001100";
WAIT FOR clk_period;
UR <= "010000010";
UI <= "000100101";
WAIT FOR clk_period;
UR <= "001111100";
UI <= "001000000";
WAIT FOR clk_period;
UR <= "001110100";
UI <= "001011100";
WAIT FOR clk_period;
UR <= "001100101";
UI <= "001110111";
WAIT FOR clk_period;
UR <= "001010001";
UI <= "010010001";
WAIT FOR clk_period;
UR <= "000110111";
UI <= "010100101";
WAIT FOR clk_period;
UR <= "000010110";
UI <= "010110001";
WAIT FOR clk_period;
UR <= "111110001";
UI <= "010111001";
WAIT FOR clk_period;
UR <= "111001001";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "110100011";
UI <= "010101101";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "010011011";
WAIT FOR clk_period;
UR <= "101100100";
UI <= "010000000";
WAIT FOR clk_period;
UR <= "101010001";
UI <= "001100000";
WAIT FOR clk_period;
UR <= "101001001";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "101001101";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "101011011";
UI <= "111101101";
WAIT FOR clk_period;
UR <= "101110010";
UI <= "111000111";
WAIT FOR clk_period;
UR <= "110010001";
UI <= "110100110";
WAIT FOR clk_period;
UR <= "110101110";
UI <= "110001011";
WAIT FOR clk_period;
UR <= "111001100";
UI <= "101110100";
WAIT FOR clk_period;
UR <= "111100000";
UI <= "101101000";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "101100010";
WAIT FOR clk_period;
UR <= "111101111";
UI <= "101100011";
WAIT FOR clk_period;
UR <= "111100100";
UI <= "101101101";
WAIT FOR clk_period;
UR <= "111001111";
UI <= "101111011";
WAIT FOR clk_period;
UR <= "110110001";
UI <= "110001111";
WAIT FOR clk_period;
UR <= "110001111";
UI <= "110101000";
WAIT FOR clk_period;
UR <= "101101111";
UI <= "111000011";
WAIT FOR clk_period;
UR <= "101010010";
UI <= "111011101";
WAIT FOR clk_period;
UR <= "100111111";
UI <= "111111000";
WAIT FOR clk_period;
UR <= "100111010";
UI <= "000010001";
WAIT FOR clk_period;
UR <= "101000110";
UI <= "000100111";
WAIT FOR clk_period;
UR <= "101100010";
UI <= "000111001";
WAIT FOR clk_period;
UR <= "110001011";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "111000000";
UI <= "001001010";
WAIT FOR clk_period;
UR <= "111111011";
UI <= "001001000";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "000101011";
WAIT FOR clk_period;
UR <= "010010111";
UI <= "000001111";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "111110001";
WAIT FOR clk_period;
UR <= "011000010";
UI <= "111001011";
WAIT FOR clk_period;
UR <= "010111110";
UI <= "110100101";
WAIT FOR clk_period;
UR <= "010101000";
UI <= "101111111";
WAIT FOR clk_period;
UR <= "010001000";
UI <= "101100000";
WAIT FOR clk_period;
UR <= "001011101";
UI <= "101001000";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "100110111";
WAIT FOR clk_period;
UR <= "000000000";
UI <= "100110010";
WAIT FOR clk_period;
UR <= "111011010";
UI <= "100111010";
WAIT FOR clk_period;
UR <= "110111100";
UI <= "101010000";
WAIT FOR clk_period;
UR <= "110101100";
UI <= "101110001";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "110011010";
WAIT FOR clk_period;
UR <= "110101111";
UI <= "111001100";
WAIT FOR clk_period;
UR <= "111000011";
UI <= "111111110";
WAIT FOR clk_period;
UR <= "111011100";
UI <= "000110001";
WAIT FOR clk_period;
UR <= "111111010";
UI <= "001011110";
WAIT FOR clk_period;
UR <= "000011000";
UI <= "010000100";
WAIT FOR clk_period;
UR <= "000110001";
UI <= "010011110";
WAIT FOR clk_period;
UR <= "001001000";
UI <= "010101100";
WAIT FOR clk_period;
UR <= "001011001";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "001100010";
UI <= "010100001";
WAIT FOR clk_period;
UR <= "001101000";
UI <= "010001010";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "001101011";
WAIT FOR clk_period;
UR <= "001101011";
UI <= "001000110";
WAIT FOR clk_period;
UR <= "001110001";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "001111001";
UI <= "111111101";
WAIT FOR clk_period;
UR <= "010000101";
UI <= "111011011";
WAIT FOR clk_period;
UR <= "010010100";
UI <= "110111111";
WAIT FOR clk_period;
UR <= "010101000";
UI <= "110101110";
WAIT FOR clk_period;
UR <= "010111011";
UI <= "110100010";
WAIT FOR clk_period;
UR <= "011001101";
UI <= "110100000";
WAIT FOR clk_period;
UR <= "011011010";
UI <= "110100010";
WAIT FOR clk_period;
UR <= "011011111";
UI <= "110101100";
WAIT FOR clk_period;
UR <= "011011100";
UI <= "110111001";
WAIT FOR clk_period;
UR <= "011010000";
UI <= "111000111";
WAIT FOR clk_period;
UR <= "010110110";
UI <= "111010111";
WAIT FOR clk_period;
UR <= "010010011";
UI <= "111100110";
WAIT FOR clk_period;
UR <= "001100110";
UI <= "111110010";
WAIT FOR clk_period;
UR <= "000110101";
UI <= "111111110";
WAIT FOR clk_period;
UR <= "000000010";
UI <= "000001000";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "000010000";
WAIT FOR clk_period;
UR <= "110100111";
UI <= "000010111";
WAIT FOR clk_period;
UR <= "110000001";
UI <= "000011101";
WAIT FOR clk_period;
UR <= "101100110";
UI <= "000100100";
WAIT FOR clk_period;
UR <= "101010111";
UI <= "000101010";
WAIT FOR clk_period;
UR <= "101010100";
UI <= "000110010";
WAIT FOR clk_period;
UR <= "101011110";
UI <= "000111011";
WAIT FOR clk_period;
UR <= "101110001";
UI <= "001000111";
WAIT FOR clk_period;
UR <= "110001010";
UI <= "001010011";
WAIT FOR clk_period;
UR <= "110101101";
UI <= "001100000";
WAIT FOR clk_period;
UR <= "111010010";
UI <= "001110001";
WAIT FOR clk_period;
UR <= "111110110";
UI <= "010000010";
WAIT FOR clk_period;
UR <= "000011001";
UI <= "010010100";
WAIT FOR clk_period;
UR <= "000111001";
UI <= "010100110";
WAIT FOR clk_period;
UR <= "001010010";
UI <= "010110111";
WAIT FOR clk_period;
UR <= "001100110";
UI <= "011000110";
WAIT FOR clk_period;
UR <= "001110001";
UI <= "011010011";
WAIT FOR clk_period;
UR <= "001110100";
UI <= "011011001";
WAIT FOR clk_period;
UR <= "001101110";
UI <= "011011010";
WAIT FOR clk_period;
UR <= "001100000";
UI <= "011010100";
WAIT FOR clk_period;
UR <= "001001100";
UI <= "011000101";
WAIT FOR clk_period;
UR <= "000110100";
UI <= "010101110";
WAIT FOR clk_period;
UR <= "000011001";
UI <= "010010000";
WAIT FOR clk_period;
UR <= "111111101";
UI <= "001101001";
WAIT FOR clk_period;
UR <= "111100011";
UI <= "000111101";
WAIT FOR clk_period;
UR <= "111001110";
UI <= "000001111";
WAIT FOR clk_period;
UR <= "110111111";
UI <= "111100000";
WAIT FOR clk_period;
UR <= "110110110";
UI <= "110110010";
WAIT FOR clk_period;
UR <= "110111000";
UI <= "110001100";
WAIT FOR clk_period;
UR <= "111000010";
UI <= "101101100";
WAIT FOR clk_period;
UR <= "111010101";
UI <= "101010111";
WAIT FOR clk_period;
UR <= "111101101";
UI <= "101001011";
WAIT FOR clk_period;
UR <= "000001011";
UI <= "101001000";
WAIT FOR clk_period;
UR <= "000101101";
UI <= "101010011";
WAIT FOR clk_period;
UR <= "001001111";
UI <= "101100011";
WAIT FOR clk_period;
UR <= "001101100";
UI <= "101111011";
WAIT FOR clk_period;
UR <= "010000101";
UI <= "110010111";
WAIT FOR clk_period;
UR <= "010011000";
UI <= "110110100";
WAIT FOR clk_period;
UR <= "010011110";
UI <= "111001111";
WAIT FOR clk_period;
UR <= "010011101";
UI <= "111100111";
WAIT FOR clk_period;
UR <= "010010001";
UI <= "111111100";
WAIT FOR clk_period;
UR <= "001111010";
UI <= "000001011";
WAIT FOR clk_period;
UR <= "001011011";
UI <= "000010110";
WAIT FOR clk_period;
UR <= "000110010";
UI <= "000011100";
WAIT FOR clk_period;
UR <= "000001000";
UI <= "000011111";
WAIT FOR clk_period;
UR <= "111011000";
UI <= "000011111";
WAIT FOR clk_period;
UR <= "110100110";
UI <= "000100000";
WAIT FOR clk_period;
UR <= "101110101";
UI <= "000100001";
WAIT FOR clk_period;
UR <= "101001010";
UI <= "000100010";
WAIT FOR clk_period;
UR <= "100100010";
UI <= "000100110";
WAIT FOR clk_period;
UR <= "100000011";
UI <= "000101011";
WAIT FOR clk_period;

      wait;
   end process;
    
END;
